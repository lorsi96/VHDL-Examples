library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sine_generator is
    port(
      clk: in std_logic;
      mul: in unsigned(3 downto 0);
      result: out std_logic
    );
end sine_generator;

architecture sine_generator_arch of sine_generator is
    signal count_ref: unsigned(7 downto 0) := "00000000";
begin
    process(clk) is
        variable address: unsigned(7 downto 0) := "00000000";
        variable counter: unsigned(8 downto 0) := "000000000";
        variable res_tmp: std_logic := '0';

    begin
        if clk = '1' then
            -- Sine Cyclic Counter --   
            if counter = count_ref then
                if counter = "11111111" then
                    res_tmp := '1';
                else
                    res_tmp := '0';
                end if;
            end if;            
            
            result <= res_tmp;

            counter := counter + 1;
            if counter = "100000000" then
                counter := "000000000";
                address := address + mul;
                if count_ref = "00000000" then
                    res_tmp := '0';
                else
                    res_tmp := '1';
                end if;
            end if;

            -- Sine Memory Map --
            case address is
                when "00000000" => count_ref <= "10000000";
                when "00000001" => count_ref <= "10000011";
                when "00000010" => count_ref <= "10000110";
                when "00000011" => count_ref <= "10001001";
                when "00000100" => count_ref <= "10001100";
                when "00000101" => count_ref <= "10001111";
                when "00000110" => count_ref <= "10010010";
                when "00000111" => count_ref <= "10010101";
                when "00001000" => count_ref <= "10011000";
                when "00001001" => count_ref <= "10011100";
                when "00001010" => count_ref <= "10011111";
                when "00001011" => count_ref <= "10100010";
                when "00001100" => count_ref <= "10100101";
                when "00001101" => count_ref <= "10101000";
                when "00001110" => count_ref <= "10101011";
                when "00001111" => count_ref <= "10101110";
                when "00010000" => count_ref <= "10110000";
                when "00010001" => count_ref <= "10110011";
                when "00010010" => count_ref <= "10110110";
                when "00010011" => count_ref <= "10111001";
                when "00010100" => count_ref <= "10111100";
                when "00010101" => count_ref <= "10111111";
                when "00010110" => count_ref <= "11000001";
                when "00010111" => count_ref <= "11000100";
                when "00011000" => count_ref <= "11000111";
                when "00011001" => count_ref <= "11001001";
                when "00011010" => count_ref <= "11001100";
                when "00011011" => count_ref <= "11001110";
                when "00011100" => count_ref <= "11010001";
                when "00011101" => count_ref <= "11010011";
                when "00011110" => count_ref <= "11010101";
                when "00011111" => count_ref <= "11011000";
                when "00100000" => count_ref <= "11011010";
                when "00100001" => count_ref <= "11011100";
                when "00100010" => count_ref <= "11011110";
                when "00100011" => count_ref <= "11100000";
                when "00100100" => count_ref <= "11100010";
                when "00100101" => count_ref <= "11100100";
                when "00100110" => count_ref <= "11100110";
                when "00100111" => count_ref <= "11101000";
                when "00101000" => count_ref <= "11101010";
                when "00101001" => count_ref <= "11101011";
                when "00101010" => count_ref <= "11101101";
                when "00101011" => count_ref <= "11101111";
                when "00101100" => count_ref <= "11110000";
                when "00101101" => count_ref <= "11110010";
                when "00101110" => count_ref <= "11110011";
                when "00101111" => count_ref <= "11110100";
                when "00110000" => count_ref <= "11110110";
                when "00110001" => count_ref <= "11110111";
                when "00110010" => count_ref <= "11111000";
                when "00110011" => count_ref <= "11111001";
                when "00110100" => count_ref <= "11111010";
                when "00110101" => count_ref <= "11111011";
                when "00110110" => count_ref <= "11111011";
                when "00110111" => count_ref <= "11111100";
                when "00111000" => count_ref <= "11111101";
                when "00111001" => count_ref <= "11111101";
                when "00111010" => count_ref <= "11111110";
                when "00111011" => count_ref <= "11111110";
                when "00111100" => count_ref <= "11111110";
                when "00111101" => count_ref <= "11111111";
                when "00111110" => count_ref <= "11111111";
                when "00111111" => count_ref <= "11111111";
                when "01000000" => count_ref <= "11111111";
                when "01000001" => count_ref <= "11111111";
                when "01000010" => count_ref <= "11111111";
                when "01000011" => count_ref <= "11111111";
                when "01000100" => count_ref <= "11111110";
                when "01000101" => count_ref <= "11111110";
                when "01000110" => count_ref <= "11111101";
                when "01000111" => count_ref <= "11111101";
                when "01001000" => count_ref <= "11111100";
                when "01001001" => count_ref <= "11111100";
                when "01001010" => count_ref <= "11111011";
                when "01001011" => count_ref <= "11111010";
                when "01001100" => count_ref <= "11111001";
                when "01001101" => count_ref <= "11111000";
                when "01001110" => count_ref <= "11110111";
                when "01001111" => count_ref <= "11110110";
                when "01010000" => count_ref <= "11110101";
                when "01010001" => count_ref <= "11110100";
                when "01010010" => count_ref <= "11110010";
                when "01010011" => count_ref <= "11110001";
                when "01010100" => count_ref <= "11101111";
                when "01010101" => count_ref <= "11101110";
                when "01010110" => count_ref <= "11101100";
                when "01010111" => count_ref <= "11101011";
                when "01011000" => count_ref <= "11101001";
                when "01011001" => count_ref <= "11100111";
                when "01011010" => count_ref <= "11100101";
                when "01011011" => count_ref <= "11100011";
                when "01011100" => count_ref <= "11100001";
                when "01011101" => count_ref <= "11011111";
                when "01011110" => count_ref <= "11011101";
                when "01011111" => count_ref <= "11011011";
                when "01100000" => count_ref <= "11011001";
                when "01100001" => count_ref <= "11010111";
                when "01100010" => count_ref <= "11010100";
                when "01100011" => count_ref <= "11010010";
                when "01100100" => count_ref <= "11001111";
                when "01100101" => count_ref <= "11001101";
                when "01100110" => count_ref <= "11001010";
                when "01100111" => count_ref <= "11001000";
                when "01101000" => count_ref <= "11000101";
                when "01101001" => count_ref <= "11000011";
                when "01101010" => count_ref <= "11000000";
                when "01101011" => count_ref <= "10111101";
                when "01101100" => count_ref <= "10111010";
                when "01101101" => count_ref <= "10111000";
                when "01101110" => count_ref <= "10110101";
                when "01101111" => count_ref <= "10110010";
                when "01110000" => count_ref <= "10101111";
                when "01110001" => count_ref <= "10101100";
                when "01110010" => count_ref <= "10101001";
                when "01110011" => count_ref <= "10100110";
                when "01110100" => count_ref <= "10100011";
                when "01110101" => count_ref <= "10100000";
                when "01110110" => count_ref <= "10011101";
                when "01110111" => count_ref <= "10011010";
                when "01111000" => count_ref <= "10010111";
                when "01111001" => count_ref <= "10010100";
                when "01111010" => count_ref <= "10010001";
                when "01111011" => count_ref <= "10001110";
                when "01111100" => count_ref <= "10001010";
                when "01111101" => count_ref <= "10000111";
                when "01111110" => count_ref <= "10000100";
                when "01111111" => count_ref <= "10000001";
                when "10000000" => count_ref <= "01111110";
                when "10000001" => count_ref <= "01111011";
                when "10000010" => count_ref <= "01111000";
                when "10000011" => count_ref <= "01110101";
                when "10000100" => count_ref <= "01110001";
                when "10000101" => count_ref <= "01101110";
                when "10000110" => count_ref <= "01101011";
                when "10000111" => count_ref <= "01101000";
                when "10001000" => count_ref <= "01100101";
                when "10001001" => count_ref <= "01100010";
                when "10001010" => count_ref <= "01011111";
                when "10001011" => count_ref <= "01011100";
                when "10001100" => count_ref <= "01011001";
                when "10001101" => count_ref <= "01010110";
                when "10001110" => count_ref <= "01010011";
                when "10001111" => count_ref <= "01010000";
                when "10010000" => count_ref <= "01001101";
                when "10010001" => count_ref <= "01001010";
                when "10010010" => count_ref <= "01000111";
                when "10010011" => count_ref <= "01000101";
                when "10010100" => count_ref <= "01000010";
                when "10010101" => count_ref <= "00111111";
                when "10010110" => count_ref <= "00111100";
                when "10010111" => count_ref <= "00111010";
                when "10011000" => count_ref <= "00110111";
                when "10011001" => count_ref <= "00110101";
                when "10011010" => count_ref <= "00110010";
                when "10011011" => count_ref <= "00110000";
                when "10011100" => count_ref <= "00101101";
                when "10011101" => count_ref <= "00101011";
                when "10011110" => count_ref <= "00101000";
                when "10011111" => count_ref <= "00100110";
                when "10100000" => count_ref <= "00100100";
                when "10100001" => count_ref <= "00100010";
                when "10100010" => count_ref <= "00100000";
                when "10100011" => count_ref <= "00011110";
                when "10100100" => count_ref <= "00011100";
                when "10100101" => count_ref <= "00011010";
                when "10100110" => count_ref <= "00011000";
                when "10100111" => count_ref <= "00010110";
                when "10101000" => count_ref <= "00010100";
                when "10101001" => count_ref <= "00010011";
                when "10101010" => count_ref <= "00010001";
                when "10101011" => count_ref <= "00010000";
                when "10101100" => count_ref <= "00001110";
                when "10101101" => count_ref <= "00001101";
                when "10101110" => count_ref <= "00001011";
                when "10101111" => count_ref <= "00001010";
                when "10110000" => count_ref <= "00001001";
                when "10110001" => count_ref <= "00001000";
                when "10110010" => count_ref <= "00000111";
                when "10110011" => count_ref <= "00000110";
                when "10110100" => count_ref <= "00000101";
                when "10110101" => count_ref <= "00000100";
                when "10110110" => count_ref <= "00000011";
                when "10110111" => count_ref <= "00000011";
                when "10111000" => count_ref <= "00000010";
                when "10111001" => count_ref <= "00000010";
                when "10111010" => count_ref <= "00000001";
                when "10111011" => count_ref <= "00000001";
                when "10111100" => count_ref <= "00000000";
                when "10111101" => count_ref <= "00000000";
                when "10111110" => count_ref <= "00000000";
                when "10111111" => count_ref <= "00000000";
                when "11000000" => count_ref <= "00000000";
                when "11000001" => count_ref <= "00000000";
                when "11000010" => count_ref <= "00000000";
                when "11000011" => count_ref <= "00000001";
                when "11000100" => count_ref <= "00000001";
                when "11000101" => count_ref <= "00000001";
                when "11000110" => count_ref <= "00000010";
                when "11000111" => count_ref <= "00000010";
                when "11001000" => count_ref <= "00000011";
                when "11001001" => count_ref <= "00000100";
                when "11001010" => count_ref <= "00000100";
                when "11001011" => count_ref <= "00000101";
                when "11001100" => count_ref <= "00000110";
                when "11001101" => count_ref <= "00000111";
                when "11001110" => count_ref <= "00001000";
                when "11001111" => count_ref <= "00001001";
                when "11010000" => count_ref <= "00001011";
                when "11010001" => count_ref <= "00001100";
                when "11010010" => count_ref <= "00001101";
                when "11010011" => count_ref <= "00001111";
                when "11010100" => count_ref <= "00010000";
                when "11010101" => count_ref <= "00010010";
                when "11010110" => count_ref <= "00010100";
                when "11010111" => count_ref <= "00010101";
                when "11011000" => count_ref <= "00010111";
                when "11011001" => count_ref <= "00011001";
                when "11011010" => count_ref <= "00011011";
                when "11011011" => count_ref <= "00011101";
                when "11011100" => count_ref <= "00011111";
                when "11011101" => count_ref <= "00100001";
                when "11011110" => count_ref <= "00100011";
                when "11011111" => count_ref <= "00100101";
                when "11100000" => count_ref <= "00100111";
                when "11100001" => count_ref <= "00101010";
                when "11100010" => count_ref <= "00101100";
                when "11100011" => count_ref <= "00101110";
                when "11100100" => count_ref <= "00110001";
                when "11100101" => count_ref <= "00110011";
                when "11100110" => count_ref <= "00110110";
                when "11100111" => count_ref <= "00111000";
                when "11101000" => count_ref <= "00111011";
                when "11101001" => count_ref <= "00111110";
                when "11101010" => count_ref <= "01000000";
                when "11101011" => count_ref <= "01000011";
                when "11101100" => count_ref <= "01000110";
                when "11101101" => count_ref <= "01001001";
                when "11101110" => count_ref <= "01001100";
                when "11101111" => count_ref <= "01001111";
                when "11110000" => count_ref <= "01010001";
                when "11110001" => count_ref <= "01010100";
                when "11110010" => count_ref <= "01010111";
                when "11110011" => count_ref <= "01011010";
                when "11110100" => count_ref <= "01011101";
                when "11110101" => count_ref <= "01100000";
                when "11110110" => count_ref <= "01100011";
                when "11110111" => count_ref <= "01100111";
                when "11111000" => count_ref <= "01101010";
                when "11111001" => count_ref <= "01101101";
                when "11111010" => count_ref <= "01110000";
                when "11111011" => count_ref <= "01110011";
                when "11111100" => count_ref <= "01110110";
                when "11111101" => count_ref <= "01111001";
                when "11111110" => count_ref <= "01111100";
                when "11111111" => count_ref <= "01111111";
                when others => count_ref <= (others => '0');
            end case;
            
        end if;
    end process;
end sine_generator_arch;   