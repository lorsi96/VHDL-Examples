library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sine_generator is
    port(
      clk: in std_logic;
      result: out std_logic_vector(7 downto 0)
    );
end sine_generator;

architecture sine_generator_arch of sine_generator is
begin
    process(clk) is
        variable address: unsigned(7 downto 0) := "00000000";
    begin
        if clk = '1' then
            -- Sine Cyclic Counter --
            -- Note: intentionally lets the counter overflow. --  
            address := address + 1;
            
            -- Sine Memory Map --
            case address is
                when "00000000" => result <= "10000000";
                when "00000001" => result <= "10000011";
                when "00000010" => result <= "10000110";
                when "00000011" => result <= "10001001";
                when "00000100" => result <= "10001100";
                when "00000101" => result <= "10001111";
                when "00000110" => result <= "10010010";
                when "00000111" => result <= "10010101";
                when "00001000" => result <= "10011000";
                when "00001001" => result <= "10011100";
                when "00001010" => result <= "10011111";
                when "00001011" => result <= "10100010";
                when "00001100" => result <= "10100101";
                when "00001101" => result <= "10101000";
                when "00001110" => result <= "10101011";
                when "00001111" => result <= "10101110";
                when "00010000" => result <= "10110000";
                when "00010001" => result <= "10110011";
                when "00010010" => result <= "10110110";
                when "00010011" => result <= "10111001";
                when "00010100" => result <= "10111100";
                when "00010101" => result <= "10111111";
                when "00010110" => result <= "11000001";
                when "00010111" => result <= "11000100";
                when "00011000" => result <= "11000111";
                when "00011001" => result <= "11001001";
                when "00011010" => result <= "11001100";
                when "00011011" => result <= "11001110";
                when "00011100" => result <= "11010001";
                when "00011101" => result <= "11010011";
                when "00011110" => result <= "11010101";
                when "00011111" => result <= "11011000";
                when "00100000" => result <= "11011010";
                when "00100001" => result <= "11011100";
                when "00100010" => result <= "11011110";
                when "00100011" => result <= "11100000";
                when "00100100" => result <= "11100010";
                when "00100101" => result <= "11100100";
                when "00100110" => result <= "11100110";
                when "00100111" => result <= "11101000";
                when "00101000" => result <= "11101010";
                when "00101001" => result <= "11101011";
                when "00101010" => result <= "11101101";
                when "00101011" => result <= "11101111";
                when "00101100" => result <= "11110000";
                when "00101101" => result <= "11110010";
                when "00101110" => result <= "11110011";
                when "00101111" => result <= "11110100";
                when "00110000" => result <= "11110110";
                when "00110001" => result <= "11110111";
                when "00110010" => result <= "11111000";
                when "00110011" => result <= "11111001";
                when "00110100" => result <= "11111010";
                when "00110101" => result <= "11111011";
                when "00110110" => result <= "11111011";
                when "00110111" => result <= "11111100";
                when "00111000" => result <= "11111101";
                when "00111001" => result <= "11111101";
                when "00111010" => result <= "11111110";
                when "00111011" => result <= "11111110";
                when "00111100" => result <= "11111110";
                when "00111101" => result <= "11111111";
                when "00111110" => result <= "11111111";
                when "00111111" => result <= "11111111";
                when "01000000" => result <= "11111111";
                when "01000001" => result <= "11111111";
                when "01000010" => result <= "11111111";
                when "01000011" => result <= "11111111";
                when "01000100" => result <= "11111110";
                when "01000101" => result <= "11111110";
                when "01000110" => result <= "11111101";
                when "01000111" => result <= "11111101";
                when "01001000" => result <= "11111100";
                when "01001001" => result <= "11111100";
                when "01001010" => result <= "11111011";
                when "01001011" => result <= "11111010";
                when "01001100" => result <= "11111001";
                when "01001101" => result <= "11111000";
                when "01001110" => result <= "11110111";
                when "01001111" => result <= "11110110";
                when "01010000" => result <= "11110101";
                when "01010001" => result <= "11110100";
                when "01010010" => result <= "11110010";
                when "01010011" => result <= "11110001";
                when "01010100" => result <= "11101111";
                when "01010101" => result <= "11101110";
                when "01010110" => result <= "11101100";
                when "01010111" => result <= "11101011";
                when "01011000" => result <= "11101001";
                when "01011001" => result <= "11100111";
                when "01011010" => result <= "11100101";
                when "01011011" => result <= "11100011";
                when "01011100" => result <= "11100001";
                when "01011101" => result <= "11011111";
                when "01011110" => result <= "11011101";
                when "01011111" => result <= "11011011";
                when "01100000" => result <= "11011001";
                when "01100001" => result <= "11010111";
                when "01100010" => result <= "11010100";
                when "01100011" => result <= "11010010";
                when "01100100" => result <= "11001111";
                when "01100101" => result <= "11001101";
                when "01100110" => result <= "11001010";
                when "01100111" => result <= "11001000";
                when "01101000" => result <= "11000101";
                when "01101001" => result <= "11000011";
                when "01101010" => result <= "11000000";
                when "01101011" => result <= "10111101";
                when "01101100" => result <= "10111010";
                when "01101101" => result <= "10111000";
                when "01101110" => result <= "10110101";
                when "01101111" => result <= "10110010";
                when "01110000" => result <= "10101111";
                when "01110001" => result <= "10101100";
                when "01110010" => result <= "10101001";
                when "01110011" => result <= "10100110";
                when "01110100" => result <= "10100011";
                when "01110101" => result <= "10100000";
                when "01110110" => result <= "10011101";
                when "01110111" => result <= "10011010";
                when "01111000" => result <= "10010111";
                when "01111001" => result <= "10010100";
                when "01111010" => result <= "10010001";
                when "01111011" => result <= "10001110";
                when "01111100" => result <= "10001010";
                when "01111101" => result <= "10000111";
                when "01111110" => result <= "10000100";
                when "01111111" => result <= "10000001";
                when "10000000" => result <= "01111110";
                when "10000001" => result <= "01111011";
                when "10000010" => result <= "01111000";
                when "10000011" => result <= "01110101";
                when "10000100" => result <= "01110001";
                when "10000101" => result <= "01101110";
                when "10000110" => result <= "01101011";
                when "10000111" => result <= "01101000";
                when "10001000" => result <= "01100101";
                when "10001001" => result <= "01100010";
                when "10001010" => result <= "01011111";
                when "10001011" => result <= "01011100";
                when "10001100" => result <= "01011001";
                when "10001101" => result <= "01010110";
                when "10001110" => result <= "01010011";
                when "10001111" => result <= "01010000";
                when "10010000" => result <= "01001101";
                when "10010001" => result <= "01001010";
                when "10010010" => result <= "01000111";
                when "10010011" => result <= "01000101";
                when "10010100" => result <= "01000010";
                when "10010101" => result <= "00111111";
                when "10010110" => result <= "00111100";
                when "10010111" => result <= "00111010";
                when "10011000" => result <= "00110111";
                when "10011001" => result <= "00110101";
                when "10011010" => result <= "00110010";
                when "10011011" => result <= "00110000";
                when "10011100" => result <= "00101101";
                when "10011101" => result <= "00101011";
                when "10011110" => result <= "00101000";
                when "10011111" => result <= "00100110";
                when "10100000" => result <= "00100100";
                when "10100001" => result <= "00100010";
                when "10100010" => result <= "00100000";
                when "10100011" => result <= "00011110";
                when "10100100" => result <= "00011100";
                when "10100101" => result <= "00011010";
                when "10100110" => result <= "00011000";
                when "10100111" => result <= "00010110";
                when "10101000" => result <= "00010100";
                when "10101001" => result <= "00010011";
                when "10101010" => result <= "00010001";
                when "10101011" => result <= "00010000";
                when "10101100" => result <= "00001110";
                when "10101101" => result <= "00001101";
                when "10101110" => result <= "00001011";
                when "10101111" => result <= "00001010";
                when "10110000" => result <= "00001001";
                when "10110001" => result <= "00001000";
                when "10110010" => result <= "00000111";
                when "10110011" => result <= "00000110";
                when "10110100" => result <= "00000101";
                when "10110101" => result <= "00000100";
                when "10110110" => result <= "00000011";
                when "10110111" => result <= "00000011";
                when "10111000" => result <= "00000010";
                when "10111001" => result <= "00000010";
                when "10111010" => result <= "00000001";
                when "10111011" => result <= "00000001";
                when "10111100" => result <= "00000000";
                when "10111101" => result <= "00000000";
                when "10111110" => result <= "00000000";
                when "10111111" => result <= "00000000";
                when "11000000" => result <= "00000000";
                when "11000001" => result <= "00000000";
                when "11000010" => result <= "00000000";
                when "11000011" => result <= "00000001";
                when "11000100" => result <= "00000001";
                when "11000101" => result <= "00000001";
                when "11000110" => result <= "00000010";
                when "11000111" => result <= "00000010";
                when "11001000" => result <= "00000011";
                when "11001001" => result <= "00000100";
                when "11001010" => result <= "00000100";
                when "11001011" => result <= "00000101";
                when "11001100" => result <= "00000110";
                when "11001101" => result <= "00000111";
                when "11001110" => result <= "00001000";
                when "11001111" => result <= "00001001";
                when "11010000" => result <= "00001011";
                when "11010001" => result <= "00001100";
                when "11010010" => result <= "00001101";
                when "11010011" => result <= "00001111";
                when "11010100" => result <= "00010000";
                when "11010101" => result <= "00010010";
                when "11010110" => result <= "00010100";
                when "11010111" => result <= "00010101";
                when "11011000" => result <= "00010111";
                when "11011001" => result <= "00011001";
                when "11011010" => result <= "00011011";
                when "11011011" => result <= "00011101";
                when "11011100" => result <= "00011111";
                when "11011101" => result <= "00100001";
                when "11011110" => result <= "00100011";
                when "11011111" => result <= "00100101";
                when "11100000" => result <= "00100111";
                when "11100001" => result <= "00101010";
                when "11100010" => result <= "00101100";
                when "11100011" => result <= "00101110";
                when "11100100" => result <= "00110001";
                when "11100101" => result <= "00110011";
                when "11100110" => result <= "00110110";
                when "11100111" => result <= "00111000";
                when "11101000" => result <= "00111011";
                when "11101001" => result <= "00111110";
                when "11101010" => result <= "01000000";
                when "11101011" => result <= "01000011";
                when "11101100" => result <= "01000110";
                when "11101101" => result <= "01001001";
                when "11101110" => result <= "01001100";
                when "11101111" => result <= "01001111";
                when "11110000" => result <= "01010001";
                when "11110001" => result <= "01010100";
                when "11110010" => result <= "01010111";
                when "11110011" => result <= "01011010";
                when "11110100" => result <= "01011101";
                when "11110101" => result <= "01100000";
                when "11110110" => result <= "01100011";
                when "11110111" => result <= "01100111";
                when "11111000" => result <= "01101010";
                when "11111001" => result <= "01101101";
                when "11111010" => result <= "01110000";
                when "11111011" => result <= "01110011";
                when "11111100" => result <= "01110110";
                when "11111101" => result <= "01111001";
                when "11111110" => result <= "01111100";
                when "11111111" => result <= "01111111";
                when others => result <= (others => 'X');
            end case;
          end if;
    end process;
end sine_generator_arch;   